module test(input x, 
				output y);
	assign y = x;
endmodule